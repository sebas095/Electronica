library ieee;use ieee.std_logic_1164.all;entity vga_test is    port(        clk     : in  std_logic;        rgb_in  : in  std_logic_vector (2 downto 0);        hsync   : out std_logic;        vsync   : out std_logic;        rgb_out : out std_logic_vector (2 downto 0)    );end vga_test;architecture Behavioral of vga_test is     component DivFreq        port(            clk  : in  std_logic;            clkout : out std_logic        );    end component;    component vga_sync        port(            pixel_clk : in  std_logic;            hsync     : out std_logic;            vsync     : out std_logic;            disp_ena  : out std_logic;            pixel_x   : out integer;            pixel_y   : out integer        );    end component;    component vga_rgb        port (            rgb_in   : in  std_logic_vector (2 downto 0);            disp_ena : in  std_logic;            rgb_out  : out std_logic_vector (2 downto 0)        );    end component;     signal pixel_clk : std_logic := '0';    signal s_disp_ena : std_logic;    signal s_pixel_x : integer;    signal s_pixel_y : integer;begin    VGA_FREQ_DIV: DivFreq port map (       clk => clk,        clkout => pixel_clk    );    VGA_SYNC_INST: vga_sync port map (        pixel_clk => pixel_clk,        hsync => hsync,        vsync => vsync,        disp_ena => s_disp_ena,        pixel_x => s_pixel_x,        pixel_y => s_pixel_y    );    VGA_RGB_INST: vga_rgb port map (        rgb_in => rgb_in,        disp_ena => s_disp_ena,        rgb_out => rgb_out    );end;